// Copyright 2018 Robert Balas <balasr@student.ethz.ch>
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

// Wrapper for a CV32E40S testbench, containing CV32E40S, Memory and stdout peripheral
// Contributor: Robert Balas <balasr@student.ethz.ch>
// Module renamed from riscv_wrapper to cv32e40s_tb_wrapper because (1) the
// name of the core changed, and (2) the design has a cv32e40s_wrapper module.
//
// SPDX-License-Identifier: Apache-2.0 WITH SHL-0.51

module cv32e40s_tb_wrapper
    #(parameter // Parameters used by TB
                INSTR_RDATA_WIDTH = 32,
                RAM_ADDR_WIDTH    = 20,
                BOOT_ADDR         = 'h80,
                DM_EXCEPTION      = 32'h1A11_1000,
                DM_HALTADDRESS    = 32'h1A11_0800,
                HART_ID           = 32'h0000_0000,
                IMP_PATCH_ID      = 4'h0,
                TRAP_VECTOR       = 32'h0000_0000
    )
    (input logic         clk_i,
     input logic         rst_ni,

     input logic         fetch_enable_i,
     output logic        tests_passed_o,
     output logic        tests_failed_o,
     output logic [31:0] exit_value_o,
     output logic        exit_valid_o);

    // signals connecting core to memory
    logic                         instr_req;
    logic                         instr_gnt;
    logic                         instr_gntpar;
    logic                         instr_rvalid;
    logic                         instr_rvalidpar;
    logic [31:0]                  instr_addr;
    logic [INSTR_RDATA_WIDTH-1:0] instr_rdata;

    logic                         data_req;
    logic                         data_gnt;
    logic                         data_gntpar;
    logic                         data_rvalid;
    logic                         data_rvalidpar;
    logic [31:0]                  data_addr;
    logic                         data_we;
    logic [3:0]                   data_be;
    logic [31:0]                  data_rdata;
    logic [31:0]                  data_wdata;

    // signals to debug unit
    logic                         debug_req;

    // irq signals (not used)
    logic [0:31]                  irq;
    logic [0:4]                   irq_id_in;
    logic                         irq_ack;
    logic [0:4]                   irq_id_out;
    logic                         irq_sec;


    // interrupts (only timer for now)
    assign irq_sec     = '0;

    assign instr_gntpar = ~instr_gnt;
    assign instr_rvalidpar = ~instr_rvalid;
    assign data_gntpar = ~data_gnt;
    assign data_rvalidpar = ~data_rvalid;
//    // core log reports parameter usage and illegal instructions to the logfile
//    // MIKET: commenting out as the cv32e40s RTL wrapper does this as well.
//    cv32e40s_core_log
//     #(
//          .PULP_XPULP            ( PULP_XPULP            ),
//          .PULP_CLUSTER          ( PULP_CLUSTER          ),
//          .FPU                   ( FPU                   ),
//          .PULP_ZFINX            ( PULP_ZFINX            ))
//    core_log_i(
//          .clk_i              ( cv32e40s_core_i.id_stage_i.clk              ),
//          .is_decoding_i      ( cv32e40s_core_i.id_stage_i.is_decoding_o    ),
//          .illegal_insn_dec_i ( cv32e40s_core_i.id_stage_i.illegal_insn_dec ),
//          .mhartid_i          ( cv32e40s_core_i.mhartid_i                   ),
//          .pc_id_i            ( cv32e40s_core_i.pc_id                       )
//      );

    // instantiate the core
    cv32e40s_core #(
          //.B_EXT                 ( ZBA_ZBB_ZBC_ZBS       ), Modified into rtl/cv32e40s_core.sv
          .DM_REGION_START       ( 32'h1A110000          ),
          .DM_REGION_END         ( 32'h1A111000          ),
          .LFSR0_CFG             ('{ coeffs : 32'h80000057, default_seed : 32'habbacafe }),
          .LFSR1_CFG             ('{ coeffs : 32'h80000062, default_seed : 32'hbeef1234 }),
          .LFSR2_CFG             ('{ coeffs : 32'h8000007a, default_seed : 32'ha5a5a5a5 })

          /// .B_EXT            (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_B_EXT),
          //.CLIC             (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC),
          //.CLIC_ID_WIDTH    (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_CLIC_ID_WIDTH),
          //.DBG_NUM_TRIGGERS (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DBG_NUM_TRIGGERS),
          /// .DM_REGION_END    (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_END),
          /// .DM_REGION_START  (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_DM_REGION_START),
          /// .LFSR0_CFG        (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_LFSR0_CFG),
          /// .LFSR1_CFG        (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_LFSR1_CFG),
          /// .LFSR2_CFG        (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_LFSR2_CFG),
          //.M_EXT            (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_M_EXT),
          //.PMA_CFG          (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_CFG),
          //.PMA_NUM_REGIONS  (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMA_NUM_REGIONS),
          //.PMP_GRANULARITY  (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_GRANULARITY),
          //.PMP_MSECCFG_RV   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_MSECCFG_RV),
          //.PMP_NUM_REGIONS  (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_NUM_REGIONS),
          //.PMP_PMPADDR_RV   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_PMPADDR_RV),
          //.PMP_PMPNCFG_RV   (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_PMP_PMPNCFG_RV),
          //.RV32             (uvmt_cv32e40s_base_test_pkg::CORE_PARAM_RV32)

         ) cv32e40s_core_i (
         .clk_i                  ( clk_i                 ),
         .rst_ni                 ( rst_ni                ),
         
         .scan_cg_en_i           ( '0                    ),

         .boot_addr_i            ( BOOT_ADDR             ),
         .dm_exception_addr_i    ( DM_EXCEPTION          ),
         .dm_halt_addr_i         ( DM_HALTADDRESS        ),
         .mhartid_i              ( HART_ID               ),
         .mimpid_patch_i         ( IMP_PATCH_ID          ),
         .mtvec_addr_i           ( TRAP_VECTOR           ),

         .instr_req_o            ( instr_req             ),
         .instr_gnt_i            ( instr_gnt             ),
         .instr_gntpar_i         ( instr_gntpar          ),
         .instr_rvalid_i         ( instr_rvalid          ),
         .instr_rvalidpar_i      ( instr_rvalidpar       ),
         .instr_addr_o           ( instr_addr            ),
         .instr_rdata_i          ( instr_rdata           ),
         .instr_err_i            ( 1'h0                  ),

         .data_req_o             ( data_req              ),
         .data_gnt_i             ( data_gnt              ),
         .data_gntpar_i          ( data_gntpar           ),
         .data_rvalid_i          ( data_rvalid           ),
         .data_rvalidpar_i       ( data_rvalidpar        ),
         .data_we_o              ( data_we               ),
         .data_be_o              ( data_be               ),
         .data_addr_o            ( data_addr             ),
         .data_wdata_o           ( data_wdata            ),
         .data_rdata_i           ( data_rdata            ),
         .data_err_i             ( 1'h0                  ),

         // Interrupts verified in UVM environment
         .irq_i                  ( {32{1'b0}}            ),
         //.irq_ack_o              ( irq_ack               ),
         //.irq_id_o               ( irq_id_out            ),
         .wu_wfe_i               ( 1'h0                  ),

         .clic_irq_i             ( 1'h0                  ),
         .clic_irq_id_i          ( 5'h00                 ),
         .clic_irq_level_i       ( 8'h00                 ),
         .clic_irq_priv_i        ( 2'h3                  ),
         .clic_irq_shv_i         ( 1'h0                  ),

         .debug_req_i            ( debug_req             ),

         .fetch_enable_i         ( fetch_enable_i        ),
         .core_sleep_o           ( core_sleep_o          )
       );

    // this handles read to RAM and memory mapped pseudo peripherals
    mm_ram
        #(.RAM_ADDR_WIDTH (RAM_ADDR_WIDTH),
          .INSTR_RDATA_WIDTH (INSTR_RDATA_WIDTH))
    ram_i
        (.clk_i          ( clk_i                                     ),
         .rst_ni         ( rst_ni                                    ),
         .dm_halt_addr_i ( DM_HALTADDRESS                            ),

         .instr_req_i    ( instr_req                                 ),
         .instr_addr_i   ( { {10{1'b0}},
                             instr_addr[RAM_ADDR_WIDTH-1:0]
                           }                                         ),
         .instr_rdata_o  ( instr_rdata                               ),
         .instr_rvalid_o ( instr_rvalid                              ),
         .instr_gnt_o    ( instr_gnt                                 ),

         .data_req_i     ( data_req                                  ),
         .data_addr_i    ( data_addr                                 ),
         .data_we_i      ( data_we                                   ),
         .data_be_i      ( data_be                                   ),
         .data_wdata_i   ( data_wdata                                ),
         .data_rdata_o   ( data_rdata                                ),
         .data_rvalid_o  ( data_rvalid                               ),
         .data_gnt_o     ( data_gnt                                  ),

         .irq_id_i       ( irq_id_out                                ),
         .irq_ack_i      ( irq_ack                                   ),
         .irq_o          ( irq                                       ),

         .debug_req_o    ( debug_req                                 ),

         .pc_core_id_i   ( cv32e40s_core_i.if_id_pipe.pc             ),

         .tests_passed_o ( tests_passed_o                            ),
         .tests_failed_o ( tests_failed_o                            ),
         .exit_valid_o   ( exit_valid_o                              ),
         .exit_value_o   ( exit_value_o                              ));

endmodule // cv32e40s_tb_wrapper
